class base_test extends uvm_test;

  function new(string name = "base_test", uvm_component parent = null);
    super.new(name,parent);
  endfunction

  extern virtual function void report_phase(uvm_phase phase);

  `uvm_component_utils(base_test)
endclass

function void base_test::report_phase(uvm_phase phase);
  uvm_report_server server;
  int err_num;

  super.report_phase(phase);

  server = get_report_server();
  err_num = server.get_severity_count(UVM_ERROR);

  if (err_num != 0) begin
    $display("TEST CASE FAILED");
  end
  else begin
    $display("TEST CASE PASSED");
  end
endfunction
