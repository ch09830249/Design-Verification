`include "my_transaction.sv"
class my_driver extends uvm_driver#(my_transaction);
    virtual my_if vif;
    virtual my_if vif2;
    `uvm_component_utils(my_driver)

    function new(string name = "my_driver", uvm_component parent = null);
        super.new(name, parent);
        `uvm_info("my_driver", "new is called", UVM_LOW);
    endfunction

    extern virtual task main_phase(uvm_phase phase);
    extern virtual task drive_one_pkt(my_transaction tr);

    virtual function void build_phase(uvm_phase phase);
        super.build_phase(phase);
        `uvm_info("my_driver", "build_phase is called", UVM_LOW);
        if(!uvm_config_db#(virtual my_if)::get(this, "", "vif", vif)) 
            `uvm_fatal("my_driver", "virtual interface must be set for vif!!!")
        else
            `uvm_info("my_driver", "get virtual interface vif successfully!!!", UVM_LOW)
    endfunction
endclass

task my_driver::main_phase(uvm_phase phase);
    vif.data <= 8'b0;
    vif.valid <= 1'b0;
    while(!vif.rst_n)
        @(posedge vif.clk);
    while(1) begin
        seq_item_port.get_next_item(req);       // 向 sequencer 發送 transaction 請求, driver 會 block 直到取得 transaction
        drive_one_pkt(req);                     // req 指向收到的 transaction, 將 transaction 分解並驅動 DUT
        seq_item_port.item_done();              // 向 sequencer 返回一個 transaction 完成的標示 
    end
    repeat(5) @(posedge vif.clk);
endtask

task my_driver::drive_one_pkt(my_transaction tr);
    byte unsigned data_q[];
    int data_size;
    
    data_size = tr.pack_bytes(data_q) / 8;
    `uvm_info("my_driver", "begin to drive one pkt", UVM_LOW);
    tr.print();
    repeat(5) @(posedge vif.clk);
    for ( int i = 0; i < data_size; i++ ) begin
        @(posedge vif.clk);
        vif.valid <= 1'b1;
        vif.data <= data_q[i];
    end

    @(posedge vif.clk);
    vif.valid <= 1'b0;
    `uvm_info("my_driver", "end drive one pkt", UVM_LOW);
endtask
